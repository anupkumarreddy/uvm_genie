/*****************************************************************************************
   filename: uart_pkg.sv
   author  : anup reddy
   description: This package contains uart uvc
******************************************************************************************/

`ifndef __uart_pkg__
   `define __uart_pkg__

/*****************************************************************************************
   Package decleration
******************************************************************************************/
package uart_pkg;
   import uvm_pkg::*
   `include "uvm_macros.svh"

/*****************************************************************************************
   Package contents
******************************************************************************************/

   `include "uart_config.sv"
   `include "uart_driver.sv"
   `include "uart_monitor.sv"
   `include "uart_sequencer.sv"
   `include "uart_agent.sv"
   `include "uart_env.sv"

endpackage : uart_pkg

`endif

/*****************************************************************************************
   End of file
******************************************************************************************/